/*
 Takes in main period signal from channel and outputs a sine wave from it.
 */
module sine_wave_generator(/*AUTOARG*/
                           // Outputs
                           sine,
                           // Inputs
                           period
                           );
   input  wire  [ 7:0] period;
   output logic [10:0] sine;

   // Brute force generated with Python
   // See sine_wave.py in this folder

   always_comb begin
      case(period)
        8'b00000000 : sine = 0;
        8'b00000001 : sine = 0;
        8'b00000010 : sine = 1;
        8'b00000011 : sine = 2;
        8'b00000100 : sine = 4;
        8'b00000101 : sine = 7;
        8'b00000110 : sine = 11;
        8'b00000111 : sine = 15;
        8'b00001000 : sine = 19;
        8'b00001001 : sine = 24;
        8'b00001010 : sine = 30;
        8'b00001011 : sine = 37;
        8'b00001100 : sine = 44;
        8'b00001101 : sine = 51;
        8'b00001110 : sine = 59;
        8'b00001111 : sine = 68;
        8'b00010000 : sine = 77;
        8'b00010001 : sine = 87;
        8'b00010010 : sine = 98;
        8'b00010011 : sine = 109;
        8'b00010100 : sine = 120;
        8'b00010101 : sine = 132;
        8'b00010110 : sine = 145;
        8'b00010111 : sine = 158;
        8'b00011000 : sine = 172;
        8'b00011001 : sine = 186;
        8'b00011010 : sine = 201;
        8'b00011011 : sine = 216;
        8'b00011100 : sine = 232;
        8'b00011101 : sine = 248;
        8'b00011110 : sine = 265;
        8'b00011111 : sine = 282;
        8'b00100000 : sine = 299;
        8'b00100001 : sine = 317;
        8'b00100010 : sine = 336;
        8'b00100011 : sine = 354;
        8'b00100100 : sine = 374;
        8'b00100101 : sine = 393;
        8'b00100110 : sine = 413;
        8'b00100111 : sine = 434;
        8'b00101000 : sine = 454;
        8'b00101001 : sine = 475;
        8'b00101010 : sine = 497;
        8'b00101011 : sine = 519;
        8'b00101100 : sine = 541;
        8'b00101101 : sine = 563;
        8'b00101110 : sine = 585;
        8'b00101111 : sine = 608;
        8'b00110000 : sine = 631;
        8'b00110001 : sine = 655;
        8'b00110010 : sine = 678;
        8'b00110011 : sine = 702;
        8'b00110100 : sine = 726;
        8'b00110101 : sine = 750;
        8'b00110110 : sine = 774;
        8'b00110111 : sine = 799;
        8'b00111000 : sine = 823;
        8'b00111001 : sine = 848;
        8'b00111010 : sine = 873;
        8'b00111011 : sine = 898;
        8'b00111100 : sine = 923;
        8'b00111101 : sine = 948;
        8'b00111110 : sine = 973;
        8'b00111111 : sine = 998;
        8'b01000000 : sine = 1023;
        8'b01000001 : sine = 1048;
        8'b01000010 : sine = 1073;
        8'b01000011 : sine = 1098;
        8'b01000100 : sine = 1123;
        8'b01000101 : sine = 1148;
        8'b01000110 : sine = 1173;
        8'b01000111 : sine = 1198;
        8'b01001000 : sine = 1223;
        8'b01001001 : sine = 1247;
        8'b01001010 : sine = 1272;
        8'b01001011 : sine = 1296;
        8'b01001100 : sine = 1320;
        8'b01001101 : sine = 1344;
        8'b01001110 : sine = 1368;
        8'b01001111 : sine = 1391;
        8'b01010000 : sine = 1415;
        8'b01010001 : sine = 1438;
        8'b01010010 : sine = 1461;
        8'b01010011 : sine = 1483;
        8'b01010100 : sine = 1505;
        8'b01010101 : sine = 1527;
        8'b01010110 : sine = 1549;
        8'b01010111 : sine = 1571;
        8'b01011000 : sine = 1592;
        8'b01011001 : sine = 1612;
        8'b01011010 : sine = 1633;
        8'b01011011 : sine = 1653;
        8'b01011100 : sine = 1672;
        8'b01011101 : sine = 1692;
        8'b01011110 : sine = 1710;
        8'b01011111 : sine = 1729;
        8'b01100000 : sine = 1747;
        8'b01100001 : sine = 1764;
        8'b01100010 : sine = 1781;
        8'b01100011 : sine = 1798;
        8'b01100100 : sine = 1814;
        8'b01100101 : sine = 1830;
        8'b01100110 : sine = 1845;
        8'b01100111 : sine = 1860;
        8'b01101000 : sine = 1874;
        8'b01101001 : sine = 1888;
        8'b01101010 : sine = 1901;
        8'b01101011 : sine = 1914;
        8'b01101100 : sine = 1926;
        8'b01101101 : sine = 1937;
        8'b01101110 : sine = 1948;
        8'b01101111 : sine = 1959;
        8'b01110000 : sine = 1969;
        8'b01110001 : sine = 1978;
        8'b01110010 : sine = 1987;
        8'b01110011 : sine = 1995;
        8'b01110100 : sine = 2002;
        8'b01110101 : sine = 2009;
        8'b01110110 : sine = 2016;
        8'b01110111 : sine = 2022;
        8'b01111000 : sine = 2027;
        8'b01111001 : sine = 2031;
        8'b01111010 : sine = 2035;
        8'b01111011 : sine = 2039;
        8'b01111100 : sine = 2042;
        8'b01111101 : sine = 2044;
        8'b01111110 : sine = 2045;
        8'b01111111 : sine = 2046;
        8'b10000000 : sine = 2047;
        8'b10000001 : sine = 2046;
        8'b10000010 : sine = 2045;
        8'b10000011 : sine = 2044;
        8'b10000100 : sine = 2042;
        8'b10000101 : sine = 2039;
        8'b10000110 : sine = 2035;
        8'b10000111 : sine = 2031;
        8'b10001000 : sine = 2027;
        8'b10001001 : sine = 2022;
        8'b10001010 : sine = 2016;
        8'b10001011 : sine = 2009;
        8'b10001100 : sine = 2002;
        8'b10001101 : sine = 1995;
        8'b10001110 : sine = 1987;
        8'b10001111 : sine = 1978;
        8'b10010000 : sine = 1969;
        8'b10010001 : sine = 1959;
        8'b10010010 : sine = 1948;
        8'b10010011 : sine = 1937;
        8'b10010100 : sine = 1926;
        8'b10010101 : sine = 1914;
        8'b10010110 : sine = 1901;
        8'b10010111 : sine = 1888;
        8'b10011000 : sine = 1874;
        8'b10011001 : sine = 1860;
        8'b10011010 : sine = 1845;
        8'b10011011 : sine = 1830;
        8'b10011100 : sine = 1814;
        8'b10011101 : sine = 1798;
        8'b10011110 : sine = 1781;
        8'b10011111 : sine = 1764;
        8'b10100000 : sine = 1747;
        8'b10100001 : sine = 1729;
        8'b10100010 : sine = 1710;
        8'b10100011 : sine = 1692;
        8'b10100100 : sine = 1672;
        8'b10100101 : sine = 1653;
        8'b10100110 : sine = 1633;
        8'b10100111 : sine = 1612;
        8'b10101000 : sine = 1592;
        8'b10101001 : sine = 1571;
        8'b10101010 : sine = 1549;
        8'b10101011 : sine = 1527;
        8'b10101100 : sine = 1505;
        8'b10101101 : sine = 1483;
        8'b10101110 : sine = 1461;
        8'b10101111 : sine = 1438;
        8'b10110000 : sine = 1415;
        8'b10110001 : sine = 1391;
        8'b10110010 : sine = 1368;
        8'b10110011 : sine = 1344;
        8'b10110100 : sine = 1320;
        8'b10110101 : sine = 1296;
        8'b10110110 : sine = 1272;
        8'b10110111 : sine = 1247;
        8'b10111000 : sine = 1223;
        8'b10111001 : sine = 1198;
        8'b10111010 : sine = 1173;
        8'b10111011 : sine = 1148;
        8'b10111100 : sine = 1123;
        8'b10111101 : sine = 1098;
        8'b10111110 : sine = 1073;
        8'b10111111 : sine = 1048;
        8'b11000000 : sine = 1023;
        8'b11000001 : sine = 998;
        8'b11000010 : sine = 973;
        8'b11000011 : sine = 948;
        8'b11000100 : sine = 923;
        8'b11000101 : sine = 898;
        8'b11000110 : sine = 873;
        8'b11000111 : sine = 848;
        8'b11001000 : sine = 823;
        8'b11001001 : sine = 799;
        8'b11001010 : sine = 774;
        8'b11001011 : sine = 750;
        8'b11001100 : sine = 726;
        8'b11001101 : sine = 702;
        8'b11001110 : sine = 678;
        8'b11001111 : sine = 655;
        8'b11010000 : sine = 631;
        8'b11010001 : sine = 608;
        8'b11010010 : sine = 585;
        8'b11010011 : sine = 563;
        8'b11010100 : sine = 541;
        8'b11010101 : sine = 519;
        8'b11010110 : sine = 497;
        8'b11010111 : sine = 475;
        8'b11011000 : sine = 454;
        8'b11011001 : sine = 434;
        8'b11011010 : sine = 413;
        8'b11011011 : sine = 393;
        8'b11011100 : sine = 374;
        8'b11011101 : sine = 354;
        8'b11011110 : sine = 336;
        8'b11011111 : sine = 317;
        8'b11100000 : sine = 299;
        8'b11100001 : sine = 282;
        8'b11100010 : sine = 265;
        8'b11100011 : sine = 248;
        8'b11100100 : sine = 232;
        8'b11100101 : sine = 216;
        8'b11100110 : sine = 201;
        8'b11100111 : sine = 186;
        8'b11101000 : sine = 172;
        8'b11101001 : sine = 158;
        8'b11101010 : sine = 145;
        8'b11101011 : sine = 132;
        8'b11101100 : sine = 120;
        8'b11101101 : sine = 109;
        8'b11101110 : sine = 98;
        8'b11101111 : sine = 87;
        8'b11110000 : sine = 77;
        8'b11110001 : sine = 68;
        8'b11110010 : sine = 59;
        8'b11110011 : sine = 51;
        8'b11110100 : sine = 44;
        8'b11110101 : sine = 37;
        8'b11110110 : sine = 30;
        8'b11110111 : sine = 24;
        8'b11111000 : sine = 19;
        8'b11111001 : sine = 15;
        8'b11111010 : sine = 11;
        8'b11111011 : sine = 7;
        8'b11111100 : sine = 4;
        8'b11111101 : sine = 2;
        8'b11111110 : sine = 1;
        8'b11111111 : sine = 0;
      endcase
   end
endmodule
