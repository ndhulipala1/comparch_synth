`default_nettype none
`timescale 1ns / 100ps


